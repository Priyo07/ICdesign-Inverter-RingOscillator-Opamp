magic
tech sky130A
magscale 1 2
timestamp 1729422526
<< nwell >>
rect 1080 2988 2472 2990
rect 1050 1754 2472 2988
rect 1080 1656 2472 1754
<< viali >>
rect 1422 1386 1554 1522
rect 1862 1384 1994 1524
rect 2276 1380 2408 1524
rect 2270 630 2318 712
<< metal1 >>
rect 1110 2958 1194 2964
rect 882 2888 1117 2958
rect 1187 2888 1824 2958
rect 1110 2882 1194 2888
rect 2168 2584 2552 2664
rect 2308 2492 2382 2494
rect 1974 2436 2382 2492
rect 1974 2428 2072 2436
rect 1260 2300 1318 2302
rect 1260 2256 1580 2300
rect 1260 1672 1318 2256
rect 1260 1614 1545 1672
rect 1441 1534 1545 1614
rect 2308 1536 2382 2436
rect 2472 1776 2552 2584
rect 2472 1696 2722 1776
rect 1118 1522 1338 1532
rect 1118 1386 1192 1522
rect 1326 1386 1338 1522
rect 1118 1376 1338 1386
rect 1416 1522 1560 1534
rect 1856 1524 2000 1536
rect 2270 1524 2414 1536
rect 1416 1386 1422 1522
rect 1554 1386 1560 1522
rect 1634 1386 1644 1522
rect 1776 1386 1786 1522
rect 1416 1374 1560 1386
rect 1856 1384 1862 1524
rect 1994 1384 2000 1524
rect 1856 1372 2000 1384
rect 2072 1380 2082 1524
rect 2214 1380 2224 1524
rect 2270 1380 2276 1524
rect 2408 1380 2414 1524
rect 1874 1310 1982 1372
rect 2270 1368 2414 1380
rect 1684 1234 1982 1310
rect 896 1078 1217 1168
rect 1127 969 1217 1078
rect 2379 995 2609 1061
rect 1127 879 1397 969
rect 2264 712 2324 724
rect 2264 630 2270 712
rect 2318 704 2324 712
rect 2379 704 2445 995
rect 2318 638 2445 704
rect 2318 630 2324 638
rect 2264 618 2324 630
rect 1135 363 1391 441
rect 656 81 734 216
rect 1135 81 1213 363
rect 656 3 1213 81
<< via1 >>
rect 1117 2888 1187 2958
rect 1192 1386 1326 1522
rect 1644 1386 1776 1522
rect 2082 1380 2214 1524
<< metal2 >>
rect 1110 2958 1194 2964
rect 1110 2888 1117 2958
rect 1187 2888 1194 2958
rect 1110 2882 1194 2888
rect 1117 1532 1187 2882
rect 1434 1824 1498 2090
rect 1434 1760 1762 1824
rect 1660 1532 1762 1760
rect 1117 1522 1338 1532
rect 1117 1417 1192 1522
rect 1118 1386 1192 1417
rect 1326 1386 1338 1522
rect 1118 1376 1338 1386
rect 1644 1522 1776 1532
rect 1644 1376 1776 1386
rect 2082 1524 2214 1534
rect 2082 1370 2214 1380
rect 1818 1294 1910 1298
rect 2102 1294 2194 1370
rect 1818 1202 2194 1294
rect 1818 892 1910 1202
<< metal3 >>
rect 528 2587 1655 2673
rect 528 2152 614 2587
rect 2196 2328 2477 2406
rect 2399 1307 2477 2328
rect 2399 1229 2819 1307
use NMOS_commonsourcegnd  NMOS_commonsourcegnd_0
timestamp 1729401142
transform 1 0 2764 0 1 137
box -258 -113 746 1903
use NMOS_RS  NMOS_RS_0
timestamp 1729221096
transform 1 0 1443 0 1 122
box -189 -100 867 1182
use PMOS_currentsource  PMOS_currentsource_0
timestamp 1729175322
transform 1 0 245 0 1 157
box -245 -167 863 2833
use PMOS_VIN_VIP_OUT  PMOS_VIN_VIP_OUT_0
timestamp 1729401836
transform 1 0 1377 0 1 2849
box -171 -1097 1051 137
<< labels >>
flabel via1 1250 1460 1250 1460 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel viali 1494 1450 1494 1450 0 FreeSans 480 0 0 0 VIP
port 1 nsew
flabel via1 1708 1444 1708 1444 0 FreeSans 480 0 0 0 OUT
port 2 nsew
flabel viali 1936 1454 1936 1454 0 FreeSans 480 0 0 0 GND
port 3 nsew
flabel via1 2156 1460 2156 1460 0 FreeSans 480 0 0 0 RS
port 4 nsew
flabel viali 2348 1450 2348 1450 0 FreeSans 480 0 0 0 VIN
port 5 nsew
<< end >>
