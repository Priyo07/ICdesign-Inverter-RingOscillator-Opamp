magic
tech sky130A
magscale 1 2
timestamp 1729401142
<< psubdiff >>
rect -241 1869 -181 1903
rect 669 1869 729 1903
rect -241 1843 -207 1869
rect 695 1843 729 1869
rect -241 -79 -207 -53
rect 695 -79 729 -53
rect -241 -113 -181 -79
rect 669 -113 729 -79
<< psubdiffcont >>
rect -181 1869 669 1903
rect -241 -53 -207 1843
rect 695 -53 729 1843
rect -181 -113 669 -79
<< poly >>
rect -90 1771 2 1787
rect -90 1737 -74 1771
rect -40 1737 2 1771
rect -90 1721 2 1737
rect -28 1703 2 1721
rect 496 1771 588 1787
rect 496 1737 538 1771
rect 572 1737 588 1771
rect 496 1721 588 1737
rect 496 1703 526 1721
rect 60 1420 220 1421
rect -90 1302 2 1318
rect 60 1312 437 1420
rect -90 1268 -74 1302
rect -40 1268 2 1302
rect -90 1252 2 1268
rect -28 1234 2 1252
rect 496 1301 588 1317
rect 496 1267 538 1301
rect 572 1267 588 1301
rect 496 1251 588 1267
rect 496 1231 526 1251
rect 60 839 438 948
rect -28 537 2 555
rect -90 521 2 537
rect -90 487 -74 521
rect -40 487 2 521
rect -90 471 2 487
rect 496 537 526 555
rect 496 521 588 537
rect 496 487 538 521
rect 572 487 588 521
rect 61 370 438 478
rect 496 471 588 487
rect 278 369 438 370
rect -28 68 2 86
rect -90 52 2 68
rect -90 18 -74 52
rect -40 18 2 52
rect -90 2 2 18
rect 496 68 526 86
rect 496 52 588 68
rect 496 18 538 52
rect 572 18 588 52
rect 496 2 588 18
<< polycont >>
rect -74 1737 -40 1771
rect 538 1737 572 1771
rect -74 1268 -40 1302
rect 538 1267 572 1301
rect -74 487 -40 521
rect 538 487 572 521
rect -74 18 -40 52
rect 538 18 572 52
<< locali >>
rect -241 1869 -181 1903
rect 669 1869 729 1903
rect -241 1843 -207 1869
rect 695 1843 729 1869
rect -90 1737 -74 1771
rect -40 1737 -24 1771
rect 522 1737 538 1771
rect 572 1737 588 1771
rect -74 1703 -39 1737
rect -74 1672 -40 1703
rect 537 1686 572 1737
rect -75 1302 -40 1303
rect -90 1268 -74 1302
rect -40 1268 -24 1302
rect -75 1234 -39 1268
rect 522 1267 538 1301
rect 572 1267 588 1301
rect -75 1206 -40 1234
rect 537 1211 572 1267
rect -75 521 -39 590
rect 538 555 572 595
rect 537 521 572 555
rect -90 487 -74 521
rect -40 487 -24 521
rect 522 487 538 521
rect 572 487 588 521
rect -74 114 -40 117
rect -74 52 -39 114
rect 537 52 572 118
rect -90 18 -74 52
rect -40 18 -24 52
rect 522 18 538 52
rect 572 18 588 52
rect -241 -79 -207 -53
rect 695 -79 729 -53
rect -241 -113 -181 -79
rect 669 -113 729 -79
<< viali >>
rect -74 1737 -40 1771
rect 538 1737 572 1771
rect -74 1268 -40 1302
rect 538 1267 572 1301
rect -252 838 -241 948
rect -241 838 -207 948
rect -207 838 -198 948
rect 686 838 695 948
rect 695 838 729 948
rect 729 838 740 948
rect -74 487 -40 521
rect 538 487 572 521
rect -74 18 -40 52
rect 538 18 572 52
<< metal1 >>
rect -86 1771 -28 1777
rect 526 1771 584 1777
rect -86 1737 -74 1771
rect -40 1737 -28 1771
rect -86 1731 -28 1737
rect 14 1737 185 1771
rect 526 1737 538 1771
rect 572 1737 584 1771
rect -74 1687 -39 1731
rect 14 1687 49 1737
rect 526 1731 584 1737
rect 537 1687 572 1731
rect -74 1685 49 1687
rect -74 1509 48 1685
rect 210 1511 220 1687
rect 278 1511 288 1687
rect 428 1511 438 1687
rect 496 1686 572 1687
rect 496 1511 571 1686
rect 451 1509 571 1511
rect -74 1508 42 1509
rect -86 1302 -28 1308
rect -86 1268 -74 1302
rect -40 1268 -28 1302
rect -86 1262 -28 1268
rect 526 1301 584 1307
rect 526 1267 538 1301
rect 572 1267 584 1301
rect -75 1219 -39 1262
rect 526 1261 584 1267
rect 537 1219 572 1261
rect -75 1217 63 1219
rect -75 1041 2 1217
rect 60 1041 70 1217
rect 210 1041 220 1217
rect 278 1041 288 1217
rect 450 1211 572 1219
rect 450 1041 570 1211
rect -75 1039 63 1041
rect 450 991 484 1041
rect -258 948 -192 960
rect 411 957 484 991
rect -258 838 -252 948
rect -198 924 -192 948
rect 680 948 746 960
rect -84 924 -24 930
rect -198 864 -84 924
rect -198 838 -192 864
rect -84 858 -24 864
rect 524 924 584 930
rect 680 924 686 948
rect 584 864 686 924
rect 524 858 584 864
rect -258 826 -192 838
rect 680 838 686 864
rect 740 838 746 948
rect 14 830 184 831
rect 13 797 184 830
rect 680 826 746 838
rect 13 749 48 797
rect -74 738 48 749
rect 450 747 570 749
rect -74 590 46 738
rect -75 571 46 590
rect 209 571 219 747
rect 277 571 287 747
rect 428 571 438 747
rect 496 595 570 747
rect 496 571 572 595
rect -75 527 -39 571
rect 537 527 572 571
rect -86 521 -28 527
rect -86 487 -74 521
rect -40 487 -28 521
rect -86 481 -28 487
rect 526 521 584 527
rect 526 487 538 521
rect 572 487 584 521
rect 526 481 584 487
rect -74 278 46 280
rect -74 102 2 278
rect 60 102 70 278
rect 210 102 220 278
rect 278 102 288 278
rect 450 118 570 279
rect -74 58 -39 102
rect 450 101 572 118
rect -86 52 -28 58
rect 450 52 484 101
rect 533 58 572 101
rect -86 18 -74 52
rect -40 18 -28 52
rect 409 18 484 52
rect 526 52 584 58
rect 526 18 538 52
rect 572 18 584 52
rect -86 12 -28 18
rect 526 12 584 18
<< via1 >>
rect 220 1511 278 1687
rect 438 1511 496 1687
rect 2 1041 60 1217
rect 220 1041 278 1217
rect -84 864 -24 924
rect 524 864 584 924
rect 219 571 277 747
rect 438 571 496 747
rect 2 102 60 278
rect 220 102 278 278
<< metal2 >>
rect 220 1687 278 1697
rect 220 1501 278 1511
rect 438 1687 496 1697
rect 438 1501 496 1511
rect 225 1227 273 1501
rect -3 1217 64 1227
rect -3 1031 64 1041
rect 220 1217 278 1227
rect 220 1031 278 1041
rect 225 924 273 1031
rect -90 864 -84 924
rect -24 864 524 924
rect 584 864 590 924
rect 225 757 273 864
rect 219 747 277 757
rect 219 561 277 571
rect 438 747 496 757
rect 438 561 496 571
rect 225 288 273 561
rect 2 278 60 288
rect 2 92 60 102
rect 220 278 278 288
rect 220 92 278 102
<< via2 >>
rect 438 1511 496 1687
rect -3 1041 2 1217
rect 2 1041 60 1217
rect 60 1041 64 1217
rect 438 571 496 747
rect 2 102 60 278
<< metal3 >>
rect 428 1687 506 1692
rect 428 1511 438 1687
rect 496 1511 506 1687
rect 428 1506 506 1511
rect -13 1217 74 1222
rect -13 1041 -3 1217
rect 64 1160 74 1217
rect 436 1160 498 1506
rect 64 1099 498 1160
rect 64 1041 74 1099
rect -13 1036 74 1041
rect 2 687 64 1036
rect 436 752 498 1099
rect 428 747 506 752
rect 428 687 438 747
rect 2 626 438 687
rect 2 283 64 626
rect 428 571 438 626
rect 496 571 506 747
rect 428 566 506 571
rect -8 278 70 283
rect -8 102 2 278
rect 60 102 70 278
rect -8 97 70 102
use sky130_fd_pr__nfet_01v8_5MNGEB  sky130_fd_pr__nfet_01v8_5MNGEB_0
timestamp 1729334380
transform 1 0 249 0 1 1599
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGEB  sky130_fd_pr__nfet_01v8_5MNGEB_1
timestamp 1729334380
transform 1 0 249 0 1 190
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGEB  sky130_fd_pr__nfet_01v8_5MNGEB_2
timestamp 1729334380
transform 1 0 249 0 1 659
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGEB  sky130_fd_pr__nfet_01v8_5MNGEB_3
timestamp 1729334380
transform 1 0 249 0 1 1129
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729334380
transform 1 0 -13 0 1 190
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729334380
transform 1 0 511 0 1 1599
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729334380
transform 1 0 511 0 1 1129
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729334380
transform 1 0 511 0 1 659
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1729334380
transform 1 0 511 0 1 190
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1729334380
transform 1 0 -13 0 1 1599
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1729334380
transform 1 0 -13 0 1 1129
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1729334380
transform 1 0 -13 0 1 659
box -73 -126 73 126
<< labels >>
flabel metal1 -52 1578 -52 1578 0 FreeSans 320 0 0 0 D8
port 0 nsew
flabel metal3 474 1364 474 1364 0 FreeSans 320 0 0 0 OUT
port 1 nsew
flabel metal1 -132 890 -132 890 0 FreeSans 320 0 0 0 GND
port 2 nsew
<< end >>
