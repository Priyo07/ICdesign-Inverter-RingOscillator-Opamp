magic
tech sky130A
magscale 1 2
timestamp 1729175322
<< nwell >>
rect -245 -167 863 2833
<< nsubdiff >>
rect -209 2763 -149 2797
rect 767 2763 827 2797
rect -209 2737 -175 2763
rect 793 2737 827 2763
rect -209 -97 -175 -71
rect 793 -97 827 -71
rect -209 -131 -149 -97
rect 767 -131 827 -97
<< nsubdiffcont >>
rect -149 2763 767 2797
rect -209 -71 -175 2737
rect 793 -71 827 2737
rect -149 -131 767 -97
<< poly >>
rect -55 2664 38 2682
rect -55 2630 -39 2664
rect -5 2630 38 2664
rect -55 2608 38 2630
rect 609 2663 702 2681
rect 609 2629 652 2663
rect 686 2629 702 2663
rect 609 2607 702 2629
rect -56 1969 37 1987
rect 94 1982 294 2088
rect -56 1935 -40 1969
rect -6 1935 37 1969
rect -56 1913 37 1935
rect 610 1969 703 1987
rect 610 1935 653 1969
rect 687 1935 703 1969
rect 610 1913 703 1935
rect 94 1238 554 1444
rect -56 746 37 768
rect -56 712 -40 746
rect -6 712 37 746
rect -56 694 37 712
rect 610 746 703 768
rect 610 712 653 746
rect 687 712 703 746
rect 352 594 552 700
rect 610 694 703 712
rect -57 52 36 74
rect -57 18 -41 52
rect -7 18 36 52
rect -57 0 36 18
rect 610 52 703 74
rect 610 18 653 52
rect 687 18 703 52
rect 610 0 703 18
<< polycont >>
rect -39 2630 -5 2664
rect 652 2629 686 2663
rect -40 1935 -6 1969
rect 653 1935 687 1969
rect -40 712 -6 746
rect 653 712 687 746
rect -41 18 -7 52
rect 653 18 687 52
<< locali >>
rect -209 2763 -149 2797
rect 767 2763 827 2797
rect -209 2737 -175 2763
rect 793 2737 827 2763
rect -55 2664 11 2681
rect -55 2630 -39 2664
rect -5 2630 11 2664
rect -55 2625 11 2630
rect 636 2663 702 2680
rect 636 2629 652 2663
rect 686 2629 702 2663
rect -40 2606 -3 2625
rect 636 2624 702 2629
rect -40 2570 -6 2606
rect 650 2570 687 2624
rect -56 1969 10 1986
rect -56 1935 -40 1969
rect -6 1935 10 1969
rect -56 1930 10 1935
rect 637 1969 703 1986
rect 637 1935 653 1969
rect 687 1935 703 1969
rect 637 1930 703 1935
rect -41 1911 -4 1930
rect -40 1873 -6 1911
rect 651 1858 688 1930
rect -40 770 -6 806
rect 652 770 686 806
rect -41 751 -4 770
rect 651 751 688 770
rect -56 746 10 751
rect -56 712 -40 746
rect -6 712 10 746
rect -56 695 10 712
rect 637 746 703 751
rect 637 712 653 746
rect 687 712 703 746
rect 637 695 703 712
rect -40 76 -6 112
rect 652 76 686 112
rect -42 57 -5 76
rect 651 57 688 76
rect -57 52 9 57
rect -57 18 -41 52
rect -7 18 9 52
rect -57 1 9 18
rect 637 52 703 57
rect 637 18 653 52
rect 687 18 703 52
rect 637 1 703 18
rect -209 -97 -175 -71
rect 793 -97 827 -71
rect -209 -131 -149 -97
rect 767 -131 827 -97
<< viali >>
rect 634 2797 702 2810
rect 634 2763 702 2797
rect 634 2750 702 2763
rect 306 2194 340 2570
rect 306 1500 340 1876
rect 306 806 340 1182
rect 306 112 340 488
rect -58 -97 8 -86
rect -58 -131 8 -97
rect -58 -140 8 -131
<< metal1 >>
rect 622 2810 714 2816
rect 622 2750 634 2810
rect 702 2750 714 2810
rect 622 2744 714 2750
rect -40 2582 -4 2667
rect 634 2624 702 2744
rect 44 2582 86 2584
rect 652 2582 688 2624
rect -62 2186 -52 2582
rect 6 2186 90 2582
rect 300 2570 346 2574
rect 300 2194 306 2570
rect 340 2194 346 2570
rect 300 2147 346 2194
rect 558 2186 700 2582
rect 558 2147 604 2186
rect 300 2101 604 2147
rect -41 1902 -7 1971
rect -46 1888 100 1902
rect -46 1486 36 1888
rect 92 1486 100 1888
rect -46 1478 100 1486
rect 300 1876 346 2101
rect 390 1934 606 1972
rect 300 1500 306 1876
rect 340 1500 346 1876
rect -52 796 90 1192
rect -40 712 -6 796
rect 42 748 90 796
rect 300 1182 346 1500
rect 554 1888 606 1934
rect 652 1888 687 1969
rect 554 1492 696 1888
rect 300 806 306 1182
rect 340 806 346 1182
rect 42 714 254 748
rect 300 581 346 806
rect 546 1196 692 1206
rect 546 794 552 1196
rect 608 794 692 1196
rect 546 782 692 794
rect 653 711 686 782
rect 42 535 346 581
rect 42 500 88 535
rect -50 104 92 500
rect 300 488 346 535
rect 300 112 306 488
rect 340 112 346 488
rect 300 108 346 112
rect 550 500 704 502
rect -40 56 -8 104
rect 44 102 84 104
rect 550 100 638 500
rect 696 100 706 500
rect -58 -80 8 56
rect 652 18 686 100
rect -70 -86 20 -80
rect -70 -140 -58 -86
rect 8 -140 20 -86
rect -70 -146 20 -140
<< via1 >>
rect -52 2186 6 2582
rect 36 1486 92 1888
rect 552 794 608 1196
rect 638 100 696 500
<< metal2 >>
rect -52 2582 6 2592
rect -52 2176 6 2186
rect -48 2082 0 2176
rect -48 2072 20 2082
rect -48 1988 20 1998
rect 630 2064 694 2073
rect 630 1991 694 2000
rect -48 696 0 1988
rect 36 1888 92 1898
rect 36 1476 92 1486
rect 36 1434 90 1476
rect 38 1376 90 1434
rect 38 1324 606 1376
rect 38 1320 90 1324
rect 554 1206 606 1324
rect 546 1196 608 1206
rect 546 794 552 1196
rect 546 782 608 794
rect -50 686 18 696
rect 638 678 694 1991
rect 627 618 636 678
rect 696 618 705 678
rect -50 604 18 614
rect 638 548 694 618
rect 638 500 696 548
rect 638 90 696 100
<< via2 >>
rect -48 1998 20 2072
rect 630 2000 694 2064
rect -50 614 18 686
rect 636 618 696 678
<< metal3 >>
rect -60 2074 52 2078
rect -60 2072 54 2074
rect -60 1998 -48 2072
rect 20 2069 54 2072
rect 20 2064 699 2069
rect 20 2000 630 2064
rect 694 2000 699 2064
rect 20 1998 699 2000
rect -60 1995 699 1998
rect -60 1994 52 1995
rect -58 1993 30 1994
rect -60 686 28 691
rect -60 614 -50 686
rect 18 684 28 686
rect 18 683 636 684
rect 18 678 701 683
rect 18 618 636 678
rect 696 618 701 678
rect 18 614 701 618
rect -60 609 28 614
rect 631 613 701 614
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729158073
transform 1 0 625 0 1 994
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729158073
transform 1 0 21 0 1 2382
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729158073
transform 1 0 625 0 1 2382
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729158073
transform 1 0 625 0 1 1688
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729158073
transform 1 0 21 0 1 1688
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729158073
transform 1 0 21 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729158073
transform 1 0 21 0 1 994
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729158073
transform 1 0 625 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729158073
transform 1 0 323 0 1 300
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729158073
transform 1 0 323 0 1 2382
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729158073
transform 1 0 323 0 1 1688
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729158073
transform 1 0 323 0 1 994
box -323 -300 323 300
<< labels >>
flabel metal1 662 2706 662 2706 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal1 580 1926 580 1926 0 FreeSans 800 0 0 0 D2
port 1 nsew
flabel metal2 60 1346 60 1346 0 FreeSans 800 0 0 0 D1
port 2 nsew
flabel metal2 664 1314 664 1314 0 FreeSans 800 0 0 0 D5
port 3 nsew
<< end >>
