magic
tech sky130A
magscale 1 2
timestamp 1729219470
<< nmos >>
rect -100 55 100 455
rect -100 -455 100 -55
<< ndiff >>
rect -158 443 -100 455
rect -158 67 -146 443
rect -112 67 -100 443
rect -158 55 -100 67
rect 100 443 158 455
rect 100 67 112 443
rect 146 67 158 443
rect 100 55 158 67
rect -158 -67 -100 -55
rect -158 -443 -146 -67
rect -112 -443 -100 -67
rect -158 -455 -100 -443
rect 100 -67 158 -55
rect 100 -443 112 -67
rect 146 -443 158 -67
rect 100 -455 158 -443
<< ndiffc >>
rect -146 67 -112 443
rect 112 67 146 443
rect -146 -443 -112 -67
rect 112 -443 146 -67
<< poly >>
rect -100 527 100 543
rect -100 493 -84 527
rect 84 493 100 527
rect -100 455 100 493
rect -100 17 100 55
rect -100 -17 -84 17
rect 84 -17 100 17
rect -100 -55 100 -17
rect -100 -493 100 -455
rect -100 -527 -84 -493
rect 84 -527 100 -493
rect -100 -543 100 -527
<< polycont >>
rect -84 493 84 527
rect -84 -17 84 17
rect -84 -527 84 -493
<< locali >>
rect -100 493 -84 527
rect 84 493 100 527
rect -146 443 -112 459
rect -146 51 -112 67
rect 112 443 146 459
rect 112 51 146 67
rect -100 -17 -84 17
rect 84 -17 100 17
rect -146 -67 -112 -51
rect -146 -459 -112 -443
rect 112 -67 146 -51
rect 112 -459 146 -443
rect -100 -527 -84 -493
rect 84 -527 100 -493
<< viali >>
rect -59 493 59 527
rect -146 67 -112 443
rect 112 67 146 443
rect -59 -17 59 17
rect -146 -443 -112 -67
rect 112 -443 146 -67
rect -59 -527 59 -493
<< metal1 >>
rect -71 527 71 533
rect -71 493 -59 527
rect 59 493 71 527
rect -71 487 71 493
rect -152 443 -106 455
rect -152 67 -146 443
rect -112 67 -106 443
rect -152 55 -106 67
rect 106 443 152 455
rect 106 67 112 443
rect 146 67 152 443
rect 106 55 152 67
rect -71 17 71 23
rect -71 -17 -59 17
rect 59 -17 71 17
rect -71 -23 71 -17
rect -152 -67 -106 -55
rect -152 -443 -146 -67
rect -112 -443 -106 -67
rect -152 -455 -106 -443
rect 106 -67 152 -55
rect 106 -443 112 -67
rect 146 -443 152 -67
rect 106 -455 152 -443
rect -71 -493 71 -487
rect -71 -527 -59 -493
rect 59 -527 71 -493
rect -71 -533 71 -527
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
