magic
tech sky130A
magscale 1 2
timestamp 1729240969
<< error_p >>
rect -36 145 36 151
rect -36 111 -24 145
rect -36 105 36 111
<< nwell >>
rect -144 -198 144 164
<< pmos >>
rect -50 -136 50 64
<< pdiff >>
rect -108 52 -50 64
rect -108 -124 -96 52
rect -62 -124 -50 52
rect -108 -136 -50 -124
rect 50 52 108 64
rect 50 -124 62 52
rect 96 -124 108 52
rect 50 -136 108 -124
<< pdiffc >>
rect -96 -124 -62 52
rect 62 -124 96 52
<< poly >>
rect -50 145 50 161
rect -50 111 -34 145
rect 34 111 50 145
rect -50 64 50 111
rect -50 -162 50 -136
<< polycont >>
rect -34 111 34 145
<< locali >>
rect -50 111 -34 145
rect 34 111 50 145
rect -96 52 -62 68
rect -96 -140 -62 -124
rect 62 52 96 68
rect 62 -140 96 -124
<< viali >>
rect -24 111 24 145
rect -96 -124 -62 52
rect 62 -124 96 52
<< metal1 >>
rect -36 145 36 151
rect -36 111 -24 145
rect 24 111 36 145
rect -36 105 36 111
rect -102 52 -56 64
rect -102 -124 -96 52
rect -62 -124 -56 52
rect -102 -136 -56 -124
rect 56 52 102 64
rect 56 -124 62 52
rect 96 -124 102 52
rect 56 -136 102 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
