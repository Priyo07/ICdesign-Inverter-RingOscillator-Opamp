magic
tech sky130A
magscale 1 2
timestamp 1729215262
<< nmos >>
rect -486 55 -86 455
rect 86 55 486 455
rect -486 -455 -86 -55
rect 86 -455 486 -55
<< ndiff >>
rect -544 443 -486 455
rect -544 67 -532 443
rect -498 67 -486 443
rect -544 55 -486 67
rect -86 443 -28 455
rect -86 67 -74 443
rect -40 67 -28 443
rect -86 55 -28 67
rect 28 443 86 455
rect 28 67 40 443
rect 74 67 86 443
rect 28 55 86 67
rect 486 443 544 455
rect 486 67 498 443
rect 532 67 544 443
rect 486 55 544 67
rect -544 -67 -486 -55
rect -544 -443 -532 -67
rect -498 -443 -486 -67
rect -544 -455 -486 -443
rect -86 -67 -28 -55
rect -86 -443 -74 -67
rect -40 -443 -28 -67
rect -86 -455 -28 -443
rect 28 -67 86 -55
rect 28 -443 40 -67
rect 74 -443 86 -67
rect 28 -455 86 -443
rect 486 -67 544 -55
rect 486 -443 498 -67
rect 532 -443 544 -67
rect 486 -455 544 -443
<< ndiffc >>
rect -532 67 -498 443
rect -74 67 -40 443
rect 40 67 74 443
rect 498 67 532 443
rect -532 -443 -498 -67
rect -74 -443 -40 -67
rect 40 -443 74 -67
rect 498 -443 532 -67
<< poly >>
rect -486 527 -86 543
rect -486 493 -470 527
rect -102 493 -86 527
rect -486 455 -86 493
rect 86 527 486 543
rect 86 493 102 527
rect 470 493 486 527
rect 86 455 486 493
rect -486 17 -86 55
rect -486 -17 -470 17
rect -102 -17 -86 17
rect -486 -55 -86 -17
rect 86 17 486 55
rect 86 -17 102 17
rect 470 -17 486 17
rect 86 -55 486 -17
rect -486 -493 -86 -455
rect -486 -527 -470 -493
rect -102 -527 -86 -493
rect -486 -543 -86 -527
rect 86 -493 486 -455
rect 86 -527 102 -493
rect 470 -527 486 -493
rect 86 -543 486 -527
<< polycont >>
rect -470 493 -102 527
rect 102 493 470 527
rect -470 -17 -102 17
rect 102 -17 470 17
rect -470 -527 -102 -493
rect 102 -527 470 -493
<< locali >>
rect -486 493 -470 527
rect -102 493 -86 527
rect 86 493 102 527
rect 470 493 486 527
rect -532 443 -498 459
rect -532 51 -498 67
rect -74 443 -40 459
rect -74 51 -40 67
rect 40 443 74 459
rect 40 51 74 67
rect 498 443 532 459
rect 498 51 532 67
rect -486 -17 -470 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 470 -17 486 17
rect -532 -67 -498 -51
rect -532 -459 -498 -443
rect -74 -67 -40 -51
rect -74 -459 -40 -443
rect 40 -67 74 -51
rect 40 -459 74 -443
rect 498 -67 532 -51
rect 498 -459 532 -443
rect -486 -527 -470 -493
rect -102 -527 -86 -493
rect 86 -527 102 -493
rect 470 -527 486 -493
<< viali >>
rect -470 493 -102 527
rect 102 493 470 527
rect -532 67 -498 443
rect -74 67 -40 443
rect 40 67 74 443
rect 498 67 532 443
rect -470 -17 -102 17
rect 102 -17 470 17
rect -532 -443 -498 -67
rect -74 -443 -40 -67
rect 40 -443 74 -67
rect 498 -443 532 -67
rect -470 -527 -102 -493
rect 102 -527 470 -493
<< metal1 >>
rect -482 527 -90 533
rect -482 493 -470 527
rect -102 493 -90 527
rect -482 487 -90 493
rect 90 527 482 533
rect 90 493 102 527
rect 470 493 482 527
rect 90 487 482 493
rect -538 443 -492 455
rect -538 67 -532 443
rect -498 67 -492 443
rect -538 55 -492 67
rect -80 443 -34 455
rect -80 67 -74 443
rect -40 67 -34 443
rect -80 55 -34 67
rect 34 443 80 455
rect 34 67 40 443
rect 74 67 80 443
rect 34 55 80 67
rect 492 443 538 455
rect 492 67 498 443
rect 532 67 538 443
rect 492 55 538 67
rect -482 17 -90 23
rect -482 -17 -470 17
rect -102 -17 -90 17
rect -482 -23 -90 -17
rect 90 17 482 23
rect 90 -17 102 17
rect 470 -17 482 17
rect 90 -23 482 -17
rect -538 -67 -492 -55
rect -538 -443 -532 -67
rect -498 -443 -492 -67
rect -538 -455 -492 -443
rect -80 -67 -34 -55
rect -80 -443 -74 -67
rect -40 -443 -34 -67
rect -80 -455 -34 -443
rect 34 -67 80 -55
rect 34 -443 40 -67
rect 74 -443 80 -67
rect 34 -455 80 -443
rect 492 -67 538 -55
rect 492 -443 498 -67
rect 532 -443 538 -67
rect 492 -455 538 -443
rect -482 -493 -90 -487
rect -482 -527 -470 -493
rect -102 -527 -90 -493
rect -482 -533 -90 -527
rect 90 -493 482 -487
rect 90 -527 102 -493
rect 470 -527 482 -493
rect 90 -533 482 -527
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 2 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
