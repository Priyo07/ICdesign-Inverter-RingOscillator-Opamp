magic
tech sky130A
magscale 1 2
timestamp 1729401836
<< nwell >>
rect -171 -1097 1051 137
<< nsubdiff >>
rect -135 67 -75 101
rect 955 67 1015 101
rect -135 41 -101 67
rect 981 41 1015 67
rect -135 -1027 -101 -1001
rect 981 -1027 1015 -1001
rect -135 -1061 -75 -1027
rect 955 -1061 1015 -1027
<< nsubdiffcont >>
rect -75 67 955 101
rect -135 -1001 -101 41
rect 981 -1001 1015 41
rect -75 -1061 955 -1027
<< poly >>
rect -12 -47 80 -30
rect -12 -81 4 -47
rect 38 -81 80 -47
rect -12 -98 80 -81
rect 50 -116 80 -98
rect 770 -45 862 -28
rect 770 -79 812 -45
rect 846 -79 862 -45
rect 770 -96 862 -79
rect 770 -114 800 -96
rect 388 -424 460 -352
rect 386 -600 458 -528
rect 48 -858 78 -840
rect -14 -875 78 -858
rect -14 -909 2 -875
rect 36 -909 78 -875
rect -14 -926 78 -909
rect 768 -858 798 -840
rect 768 -875 860 -858
rect 768 -909 810 -875
rect 844 -909 860 -875
rect 768 -926 860 -909
<< polycont >>
rect 4 -81 38 -47
rect 812 -79 846 -45
rect 2 -909 36 -875
rect 810 -909 844 -875
<< locali >>
rect -135 67 -75 101
rect 955 67 1015 101
rect -135 41 -101 67
rect 981 41 1015 67
rect 4 -47 38 -46
rect -12 -81 4 -47
rect 38 -81 54 -47
rect 796 -79 812 -45
rect 846 -79 862 -45
rect 4 -154 38 -81
rect 812 -160 846 -79
rect 2 -875 36 -798
rect 810 -875 844 -790
rect -14 -909 2 -875
rect 36 -909 52 -875
rect 794 -909 810 -875
rect 844 -909 860 -875
rect 2 -910 36 -909
rect -135 -1027 -101 -1001
rect 981 -1027 1015 -1001
rect -135 -1061 -75 -1027
rect 955 -1061 1015 -1027
<< viali >>
rect 388 101 462 104
rect 388 67 462 101
rect 388 62 462 67
rect 4 -81 38 -47
rect 812 -79 846 -45
rect 2 -909 36 -875
rect 810 -909 844 -875
rect 386 -1027 460 -1024
rect 386 -1061 460 -1027
rect 386 -1066 460 -1061
<< metal1 >>
rect 376 104 474 110
rect 376 62 388 104
rect 462 62 474 104
rect 376 56 474 62
rect 390 -12 462 -4
rect -8 -47 50 -41
rect -8 -81 4 -47
rect 38 -81 50 -47
rect 390 -72 396 -12
rect 456 -18 462 -12
rect 458 -70 462 -18
rect 456 -72 462 -70
rect 390 -80 462 -72
rect 800 -45 858 -39
rect 800 -79 812 -45
rect 846 -79 858 -45
rect -8 -87 50 -81
rect 4 -138 38 -87
rect -18 -140 44 -138
rect -18 -318 128 -140
rect 232 -316 242 -140
rect 294 -316 304 -140
rect -18 -440 38 -318
rect 396 -322 456 -80
rect 800 -85 858 -79
rect 812 -140 846 -85
rect 546 -316 556 -140
rect 608 -316 618 -140
rect 704 -316 714 -140
rect 768 -316 848 -140
rect 724 -318 848 -316
rect 152 -418 162 -366
rect 214 -418 224 -366
rect 310 -416 382 -370
rect 466 -376 542 -362
rect -28 -452 50 -440
rect 321 -451 371 -416
rect 458 -418 548 -376
rect 622 -418 632 -364
rect 686 -368 696 -364
rect 686 -416 698 -368
rect 686 -418 696 -416
rect -28 -508 -18 -452
rect 38 -508 50 -452
rect -28 -520 50 -508
rect 160 -501 371 -451
rect 480 -458 528 -418
rect 824 -454 902 -442
rect 160 -540 210 -501
rect 480 -506 684 -458
rect 314 -536 372 -530
rect 150 -546 222 -540
rect 136 -586 236 -546
rect 308 -588 318 -536
rect 370 -588 380 -536
rect 466 -588 476 -534
rect 530 -588 540 -534
rect 636 -536 684 -506
rect 824 -510 834 -454
rect 890 -510 902 -454
rect 824 -524 902 -510
rect 616 -590 706 -536
rect 0 -638 124 -636
rect 0 -814 80 -638
rect 134 -814 144 -638
rect 230 -814 240 -638
rect 292 -814 302 -638
rect 2 -869 36 -814
rect -10 -875 48 -869
rect 394 -874 454 -622
rect 834 -636 890 -524
rect 544 -814 554 -638
rect 606 -814 616 -638
rect 720 -814 890 -636
rect 810 -822 890 -814
rect 810 -869 844 -822
rect -10 -909 2 -875
rect 36 -909 48 -875
rect -10 -915 48 -909
rect 386 -882 460 -874
rect 386 -942 394 -882
rect 454 -942 460 -882
rect 798 -875 856 -869
rect 798 -909 810 -875
rect 844 -909 856 -875
rect 798 -915 856 -909
rect 386 -948 460 -942
rect 374 -1024 472 -1018
rect 374 -1066 386 -1024
rect 460 -1066 472 -1024
rect 374 -1072 472 -1066
<< via1 >>
rect 396 -18 456 -12
rect 396 -70 458 -18
rect 396 -72 456 -70
rect 242 -316 294 -140
rect 556 -316 608 -140
rect 714 -316 768 -140
rect 162 -418 214 -366
rect 632 -418 686 -364
rect -18 -508 38 -452
rect 318 -588 370 -536
rect 476 -588 530 -534
rect 834 -510 890 -454
rect 80 -814 134 -638
rect 240 -814 292 -638
rect 554 -814 606 -638
rect 394 -942 454 -882
<< metal2 >>
rect 390 -12 462 -4
rect 390 -18 396 -12
rect 80 -70 396 -18
rect 456 -18 462 -12
rect 458 -70 464 -18
rect -28 -450 50 -440
rect -28 -510 -20 -450
rect 40 -510 50 -450
rect -28 -520 50 -510
rect 80 -628 132 -70
rect 390 -72 396 -70
rect 456 -72 462 -70
rect 390 -80 462 -72
rect 240 -140 296 -130
rect 240 -326 296 -316
rect 554 -140 610 -130
rect 554 -326 610 -316
rect 714 -140 768 -130
rect 714 -326 768 -316
rect 162 -366 214 -356
rect 632 -363 686 -354
rect 632 -364 687 -363
rect 214 -418 218 -368
rect 162 -450 218 -418
rect 686 -418 687 -364
rect 632 -450 687 -418
rect 162 -506 374 -450
rect 316 -536 374 -506
rect 316 -580 318 -536
rect 370 -580 374 -536
rect 476 -504 687 -450
rect 476 -534 530 -504
rect 370 -586 372 -580
rect 318 -598 370 -588
rect 476 -598 530 -588
rect 80 -638 134 -628
rect 80 -824 134 -814
rect 238 -638 294 -628
rect 238 -824 294 -814
rect 552 -638 608 -628
rect 552 -824 608 -814
rect 386 -882 460 -874
rect 386 -942 394 -882
rect 454 -891 460 -882
rect 718 -891 768 -326
rect 824 -452 902 -442
rect 824 -512 832 -452
rect 892 -512 902 -452
rect 824 -524 902 -512
rect 454 -941 768 -891
rect 454 -942 460 -941
rect 386 -948 460 -942
<< via2 >>
rect 398 -70 454 -14
rect -20 -452 40 -450
rect -20 -508 -18 -452
rect -18 -508 38 -452
rect 38 -508 40 -452
rect -20 -510 40 -508
rect 240 -316 242 -140
rect 242 -316 294 -140
rect 294 -316 296 -140
rect 554 -316 556 -140
rect 556 -316 608 -140
rect 608 -316 610 -140
rect 238 -814 240 -638
rect 240 -814 292 -638
rect 292 -814 294 -638
rect 552 -814 554 -638
rect 554 -814 606 -638
rect 606 -814 608 -638
rect 396 -940 452 -884
rect 832 -454 892 -452
rect 832 -510 834 -454
rect 834 -510 890 -454
rect 890 -510 892 -454
rect 832 -512 892 -510
<< metal3 >>
rect 390 -12 462 -4
rect 390 -14 892 -12
rect 390 -70 398 -14
rect 454 -70 892 -14
rect 390 -72 892 -70
rect 390 -80 462 -72
rect 230 -140 306 -135
rect 230 -316 240 -140
rect 296 -184 306 -140
rect 544 -140 620 -135
rect 544 -184 554 -140
rect 296 -246 554 -184
rect 296 -316 306 -246
rect 230 -321 306 -316
rect -28 -450 50 -440
rect -28 -510 -20 -450
rect 40 -510 50 -450
rect -28 -520 50 -510
rect -20 -882 40 -520
rect 228 -638 304 -633
rect 228 -814 238 -638
rect 294 -692 304 -638
rect 386 -692 462 -246
rect 544 -316 554 -246
rect 610 -316 620 -140
rect 544 -321 620 -316
rect 832 -442 892 -72
rect 824 -452 902 -442
rect 824 -512 832 -452
rect 892 -512 902 -452
rect 824 -524 902 -512
rect 542 -638 618 -633
rect 542 -692 552 -638
rect 294 -754 552 -692
rect 294 -814 304 -754
rect 228 -819 304 -814
rect 542 -814 552 -754
rect 608 -814 618 -638
rect 542 -819 618 -814
rect 386 -882 460 -874
rect -20 -884 460 -882
rect -20 -940 396 -884
rect 452 -940 460 -884
rect -20 -942 460 -940
rect 386 -948 460 -942
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729233510
transform 1 0 63 0 1 -726
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729233510
transform 1 0 65 0 1 -228
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729233510
transform 1 0 783 0 1 -726
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729233510
transform 1 0 785 0 1 -228
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_4TGZK8  sky130_fd_pr__pfet_01v8_4TGZK8_0
timestamp 1729240969
transform 1 0 660 0 1 -690
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_4TGZK8  sky130_fd_pr__pfet_01v8_4TGZK8_1
timestamp 1729240969
transform 1 0 502 0 1 -690
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_4TGZK8  sky130_fd_pr__pfet_01v8_4TGZK8_2
timestamp 1729240969
transform 1 0 344 0 1 -690
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_4TGZK8  sky130_fd_pr__pfet_01v8_4TGZK8_3
timestamp 1729240969
transform 1 0 186 0 1 -690
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_7WEZ7N  sky130_fd_pr__pfet_01v8_7WEZ7N_0
timestamp 1729235384
transform 1 0 346 0 1 -264
box -144 -164 144 198
use sky130_fd_pr__pfet_01v8_7WEZ7N  sky130_fd_pr__pfet_01v8_7WEZ7N_1
timestamp 1729235384
transform 1 0 188 0 1 -264
box -144 -164 144 198
use sky130_fd_pr__pfet_01v8_7WEZ7N  sky130_fd_pr__pfet_01v8_7WEZ7N_2
timestamp 1729235384
transform 1 0 662 0 1 -264
box -144 -164 144 198
use sky130_fd_pr__pfet_01v8_7WEZ7N  sky130_fd_pr__pfet_01v8_7WEZ7N_3
timestamp 1729235384
transform 1 0 504 0 1 -264
box -144 -164 144 198
<< labels >>
flabel metal1 190 -520 190 -520 0 FreeSans 480 0 0 0 VIP
port 0 nsew
flabel metal2 652 -438 652 -438 0 FreeSans 480 0 0 0 VIN
port 1 nsew
flabel viali 434 78 434 78 0 FreeSans 480 0 0 0 VDD
port 2 nsew
flabel metal1 4 -390 4 -390 0 FreeSans 480 0 0 0 D6
port 3 nsew
flabel metal3 860 -396 860 -396 0 FreeSans 480 0 0 0 OUT
port 4 nsew
flabel metal3 340 -218 340 -218 0 FreeSans 480 0 0 0 D5
port 5 nsew
<< end >>
